[Foo]
U32 state
U64 time
I8 a
I16 b
I32 c
I64 d
U8 e
U16 f
U32 g
U64 h
F32 i
F64 j
BOOL k
