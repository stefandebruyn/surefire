[Foo]
U32 state
U64 time
U64 n
U64 fib_n
