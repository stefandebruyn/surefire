[Foo]
U32 state
U64 time
F64 altitude
F64 verticalVelocity
bool enableEngine
bool popNosecone
bool deployParachute
bool ventOpen
