[Foo]
I32 foo
F64 bar
U32 state
U64 time

[Bar]
BOOL baz
