[Foo]
U32 state
U64 time
I8 a
I16 b
I32 c
I64 d
U8 e
U16 f
U32 g
U64 h
F32 i
F64 j
bool k
I32 foo
I32 bar
I32 baz
F64 qux
F64 corge
F64 grault
I8 alpha_sv
I16 beta_sv
I32 gamma_sv
I64 delta_sv
U8 epsilon_sv
U16 zeta_sv
U32 eta_sv
U64 theta_sv
F32 iota_sv
F64 kappa_sv
bool lambda_sv
F64 pi_sv
F64 tau_sv
F32 euler_sv
